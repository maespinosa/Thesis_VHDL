-------------------------------------------------------------------------------
--
-- Title       : Convolution_Layer_Top
-- Design      : Convolution_Layer
-- Author      : Marks-M3800
-- Company     : Cal Poly Pomona
--
-------------------------------------------------------------------------------
--
-- File        : C:\Sourcetree_Local\Thesis_VHDL\Active_HDL_Projects\Convolution_Layer\Convolution_Layer\compile\Convolution_Layer_Top.vhd
-- Generated   : Sat Aug 12 16:47:46 2017
-- From        : C:\Sourcetree_Local\Thesis_VHDL\Active_HDL_Projects\Convolution_Layer\Convolution_Layer\src\Convolution_Layer_Top.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;


entity Convolution_Layer_Top is 
end Convolution_Layer_Top;

architecture arch of Convolution_Layer_Top is

---- Component declarations -----

component Convolution_Controller
  port (
       i_clear_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_clk : in STD_LOGIC;
       i_conv_parameters_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_filter_data_addr_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_filter_data_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_input_data_addr_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_input_data_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_output_data_addr_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_output_data_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_relu_control_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_repeat_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_reset_n : in STD_LOGIC;
       i_start_reg : in STD_LOGIC_VECTOR(31 downto 0);
       i_status_reg : in STD_LOGIC_VECTOR(31 downto 0);
       o_clear_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_conv_parameters_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_filter_data_addr_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_filter_data_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_input_data_addr_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_input_data_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_output_data_addr_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_output_data_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_relu_control_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_repeat_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_start_reg : out STD_LOGIC_VECTOR(31 downto 0);
       o_status_reg : out STD_LOGIC_VECTOR(31 downto 0)
  );
end component;

----     Constants     -----
constant DANGLING_INPUT_CONSTANT : STD_LOGIC := 'Z';

---- Declaration for Dangling input ----
signal Dangling_Input_Signal : STD_LOGIC;

begin

----  Component instantiations  ----

U1 : Convolution_Controller
  port map(
       i_clear_reg(0) => Dangling_Input_Signal,
       i_clear_reg(1) => Dangling_Input_Signal,
       i_clear_reg(2) => Dangling_Input_Signal,
       i_clear_reg(3) => Dangling_Input_Signal,
       i_clear_reg(4) => Dangling_Input_Signal,
       i_clear_reg(5) => Dangling_Input_Signal,
       i_clear_reg(6) => Dangling_Input_Signal,
       i_clear_reg(7) => Dangling_Input_Signal,
       i_clear_reg(8) => Dangling_Input_Signal,
       i_clear_reg(9) => Dangling_Input_Signal,
       i_clear_reg(10) => Dangling_Input_Signal,
       i_clear_reg(11) => Dangling_Input_Signal,
       i_clear_reg(12) => Dangling_Input_Signal,
       i_clear_reg(13) => Dangling_Input_Signal,
       i_clear_reg(14) => Dangling_Input_Signal,
       i_clear_reg(15) => Dangling_Input_Signal,
       i_clear_reg(16) => Dangling_Input_Signal,
       i_clear_reg(17) => Dangling_Input_Signal,
       i_clear_reg(18) => Dangling_Input_Signal,
       i_clear_reg(19) => Dangling_Input_Signal,
       i_clear_reg(20) => Dangling_Input_Signal,
       i_clear_reg(21) => Dangling_Input_Signal,
       i_clear_reg(22) => Dangling_Input_Signal,
       i_clear_reg(23) => Dangling_Input_Signal,
       i_clear_reg(24) => Dangling_Input_Signal,
       i_clear_reg(25) => Dangling_Input_Signal,
       i_clear_reg(26) => Dangling_Input_Signal,
       i_clear_reg(27) => Dangling_Input_Signal,
       i_clear_reg(28) => Dangling_Input_Signal,
       i_clear_reg(29) => Dangling_Input_Signal,
       i_clear_reg(30) => Dangling_Input_Signal,
       i_clear_reg(31) => Dangling_Input_Signal,
       i_conv_parameters_reg(0) => Dangling_Input_Signal,
       i_conv_parameters_reg(1) => Dangling_Input_Signal,
       i_conv_parameters_reg(2) => Dangling_Input_Signal,
       i_conv_parameters_reg(3) => Dangling_Input_Signal,
       i_conv_parameters_reg(4) => Dangling_Input_Signal,
       i_conv_parameters_reg(5) => Dangling_Input_Signal,
       i_conv_parameters_reg(6) => Dangling_Input_Signal,
       i_conv_parameters_reg(7) => Dangling_Input_Signal,
       i_conv_parameters_reg(8) => Dangling_Input_Signal,
       i_conv_parameters_reg(9) => Dangling_Input_Signal,
       i_conv_parameters_reg(10) => Dangling_Input_Signal,
       i_conv_parameters_reg(11) => Dangling_Input_Signal,
       i_conv_parameters_reg(12) => Dangling_Input_Signal,
       i_conv_parameters_reg(13) => Dangling_Input_Signal,
       i_conv_parameters_reg(14) => Dangling_Input_Signal,
       i_conv_parameters_reg(15) => Dangling_Input_Signal,
       i_conv_parameters_reg(16) => Dangling_Input_Signal,
       i_conv_parameters_reg(17) => Dangling_Input_Signal,
       i_conv_parameters_reg(18) => Dangling_Input_Signal,
       i_conv_parameters_reg(19) => Dangling_Input_Signal,
       i_conv_parameters_reg(20) => Dangling_Input_Signal,
       i_conv_parameters_reg(21) => Dangling_Input_Signal,
       i_conv_parameters_reg(22) => Dangling_Input_Signal,
       i_conv_parameters_reg(23) => Dangling_Input_Signal,
       i_conv_parameters_reg(24) => Dangling_Input_Signal,
       i_conv_parameters_reg(25) => Dangling_Input_Signal,
       i_conv_parameters_reg(26) => Dangling_Input_Signal,
       i_conv_parameters_reg(27) => Dangling_Input_Signal,
       i_conv_parameters_reg(28) => Dangling_Input_Signal,
       i_conv_parameters_reg(29) => Dangling_Input_Signal,
       i_conv_parameters_reg(30) => Dangling_Input_Signal,
       i_conv_parameters_reg(31) => Dangling_Input_Signal,
       i_filter_data_addr_reg(0) => Dangling_Input_Signal,
       i_filter_data_addr_reg(1) => Dangling_Input_Signal,
       i_filter_data_addr_reg(2) => Dangling_Input_Signal,
       i_filter_data_addr_reg(3) => Dangling_Input_Signal,
       i_filter_data_addr_reg(4) => Dangling_Input_Signal,
       i_filter_data_addr_reg(5) => Dangling_Input_Signal,
       i_filter_data_addr_reg(6) => Dangling_Input_Signal,
       i_filter_data_addr_reg(7) => Dangling_Input_Signal,
       i_filter_data_addr_reg(8) => Dangling_Input_Signal,
       i_filter_data_addr_reg(9) => Dangling_Input_Signal,
       i_filter_data_addr_reg(10) => Dangling_Input_Signal,
       i_filter_data_addr_reg(11) => Dangling_Input_Signal,
       i_filter_data_addr_reg(12) => Dangling_Input_Signal,
       i_filter_data_addr_reg(13) => Dangling_Input_Signal,
       i_filter_data_addr_reg(14) => Dangling_Input_Signal,
       i_filter_data_addr_reg(15) => Dangling_Input_Signal,
       i_filter_data_addr_reg(16) => Dangling_Input_Signal,
       i_filter_data_addr_reg(17) => Dangling_Input_Signal,
       i_filter_data_addr_reg(18) => Dangling_Input_Signal,
       i_filter_data_addr_reg(19) => Dangling_Input_Signal,
       i_filter_data_addr_reg(20) => Dangling_Input_Signal,
       i_filter_data_addr_reg(21) => Dangling_Input_Signal,
       i_filter_data_addr_reg(22) => Dangling_Input_Signal,
       i_filter_data_addr_reg(23) => Dangling_Input_Signal,
       i_filter_data_addr_reg(24) => Dangling_Input_Signal,
       i_filter_data_addr_reg(25) => Dangling_Input_Signal,
       i_filter_data_addr_reg(26) => Dangling_Input_Signal,
       i_filter_data_addr_reg(27) => Dangling_Input_Signal,
       i_filter_data_addr_reg(28) => Dangling_Input_Signal,
       i_filter_data_addr_reg(29) => Dangling_Input_Signal,
       i_filter_data_addr_reg(30) => Dangling_Input_Signal,
       i_filter_data_addr_reg(31) => Dangling_Input_Signal,
       i_filter_data_reg(0) => Dangling_Input_Signal,
       i_filter_data_reg(1) => Dangling_Input_Signal,
       i_filter_data_reg(2) => Dangling_Input_Signal,
       i_filter_data_reg(3) => Dangling_Input_Signal,
       i_filter_data_reg(4) => Dangling_Input_Signal,
       i_filter_data_reg(5) => Dangling_Input_Signal,
       i_filter_data_reg(6) => Dangling_Input_Signal,
       i_filter_data_reg(7) => Dangling_Input_Signal,
       i_filter_data_reg(8) => Dangling_Input_Signal,
       i_filter_data_reg(9) => Dangling_Input_Signal,
       i_filter_data_reg(10) => Dangling_Input_Signal,
       i_filter_data_reg(11) => Dangling_Input_Signal,
       i_filter_data_reg(12) => Dangling_Input_Signal,
       i_filter_data_reg(13) => Dangling_Input_Signal,
       i_filter_data_reg(14) => Dangling_Input_Signal,
       i_filter_data_reg(15) => Dangling_Input_Signal,
       i_filter_data_reg(16) => Dangling_Input_Signal,
       i_filter_data_reg(17) => Dangling_Input_Signal,
       i_filter_data_reg(18) => Dangling_Input_Signal,
       i_filter_data_reg(19) => Dangling_Input_Signal,
       i_filter_data_reg(20) => Dangling_Input_Signal,
       i_filter_data_reg(21) => Dangling_Input_Signal,
       i_filter_data_reg(22) => Dangling_Input_Signal,
       i_filter_data_reg(23) => Dangling_Input_Signal,
       i_filter_data_reg(24) => Dangling_Input_Signal,
       i_filter_data_reg(25) => Dangling_Input_Signal,
       i_filter_data_reg(26) => Dangling_Input_Signal,
       i_filter_data_reg(27) => Dangling_Input_Signal,
       i_filter_data_reg(28) => Dangling_Input_Signal,
       i_filter_data_reg(29) => Dangling_Input_Signal,
       i_filter_data_reg(30) => Dangling_Input_Signal,
       i_filter_data_reg(31) => Dangling_Input_Signal,
       i_input_data_addr_reg(0) => Dangling_Input_Signal,
       i_input_data_addr_reg(1) => Dangling_Input_Signal,
       i_input_data_addr_reg(2) => Dangling_Input_Signal,
       i_input_data_addr_reg(3) => Dangling_Input_Signal,
       i_input_data_addr_reg(4) => Dangling_Input_Signal,
       i_input_data_addr_reg(5) => Dangling_Input_Signal,
       i_input_data_addr_reg(6) => Dangling_Input_Signal,
       i_input_data_addr_reg(7) => Dangling_Input_Signal,
       i_input_data_addr_reg(8) => Dangling_Input_Signal,
       i_input_data_addr_reg(9) => Dangling_Input_Signal,
       i_input_data_addr_reg(10) => Dangling_Input_Signal,
       i_input_data_addr_reg(11) => Dangling_Input_Signal,
       i_input_data_addr_reg(12) => Dangling_Input_Signal,
       i_input_data_addr_reg(13) => Dangling_Input_Signal,
       i_input_data_addr_reg(14) => Dangling_Input_Signal,
       i_input_data_addr_reg(15) => Dangling_Input_Signal,
       i_input_data_addr_reg(16) => Dangling_Input_Signal,
       i_input_data_addr_reg(17) => Dangling_Input_Signal,
       i_input_data_addr_reg(18) => Dangling_Input_Signal,
       i_input_data_addr_reg(19) => Dangling_Input_Signal,
       i_input_data_addr_reg(20) => Dangling_Input_Signal,
       i_input_data_addr_reg(21) => Dangling_Input_Signal,
       i_input_data_addr_reg(22) => Dangling_Input_Signal,
       i_input_data_addr_reg(23) => Dangling_Input_Signal,
       i_input_data_addr_reg(24) => Dangling_Input_Signal,
       i_input_data_addr_reg(25) => Dangling_Input_Signal,
       i_input_data_addr_reg(26) => Dangling_Input_Signal,
       i_input_data_addr_reg(27) => Dangling_Input_Signal,
       i_input_data_addr_reg(28) => Dangling_Input_Signal,
       i_input_data_addr_reg(29) => Dangling_Input_Signal,
       i_input_data_addr_reg(30) => Dangling_Input_Signal,
       i_input_data_addr_reg(31) => Dangling_Input_Signal,
       i_input_data_reg(0) => Dangling_Input_Signal,
       i_input_data_reg(1) => Dangling_Input_Signal,
       i_input_data_reg(2) => Dangling_Input_Signal,
       i_input_data_reg(3) => Dangling_Input_Signal,
       i_input_data_reg(4) => Dangling_Input_Signal,
       i_input_data_reg(5) => Dangling_Input_Signal,
       i_input_data_reg(6) => Dangling_Input_Signal,
       i_input_data_reg(7) => Dangling_Input_Signal,
       i_input_data_reg(8) => Dangling_Input_Signal,
       i_input_data_reg(9) => Dangling_Input_Signal,
       i_input_data_reg(10) => Dangling_Input_Signal,
       i_input_data_reg(11) => Dangling_Input_Signal,
       i_input_data_reg(12) => Dangling_Input_Signal,
       i_input_data_reg(13) => Dangling_Input_Signal,
       i_input_data_reg(14) => Dangling_Input_Signal,
       i_input_data_reg(15) => Dangling_Input_Signal,
       i_input_data_reg(16) => Dangling_Input_Signal,
       i_input_data_reg(17) => Dangling_Input_Signal,
       i_input_data_reg(18) => Dangling_Input_Signal,
       i_input_data_reg(19) => Dangling_Input_Signal,
       i_input_data_reg(20) => Dangling_Input_Signal,
       i_input_data_reg(21) => Dangling_Input_Signal,
       i_input_data_reg(22) => Dangling_Input_Signal,
       i_input_data_reg(23) => Dangling_Input_Signal,
       i_input_data_reg(24) => Dangling_Input_Signal,
       i_input_data_reg(25) => Dangling_Input_Signal,
       i_input_data_reg(26) => Dangling_Input_Signal,
       i_input_data_reg(27) => Dangling_Input_Signal,
       i_input_data_reg(28) => Dangling_Input_Signal,
       i_input_data_reg(29) => Dangling_Input_Signal,
       i_input_data_reg(30) => Dangling_Input_Signal,
       i_input_data_reg(31) => Dangling_Input_Signal,
       i_output_data_addr_reg(0) => Dangling_Input_Signal,
       i_output_data_addr_reg(1) => Dangling_Input_Signal,
       i_output_data_addr_reg(2) => Dangling_Input_Signal,
       i_output_data_addr_reg(3) => Dangling_Input_Signal,
       i_output_data_addr_reg(4) => Dangling_Input_Signal,
       i_output_data_addr_reg(5) => Dangling_Input_Signal,
       i_output_data_addr_reg(6) => Dangling_Input_Signal,
       i_output_data_addr_reg(7) => Dangling_Input_Signal,
       i_output_data_addr_reg(8) => Dangling_Input_Signal,
       i_output_data_addr_reg(9) => Dangling_Input_Signal,
       i_output_data_addr_reg(10) => Dangling_Input_Signal,
       i_output_data_addr_reg(11) => Dangling_Input_Signal,
       i_output_data_addr_reg(12) => Dangling_Input_Signal,
       i_output_data_addr_reg(13) => Dangling_Input_Signal,
       i_output_data_addr_reg(14) => Dangling_Input_Signal,
       i_output_data_addr_reg(15) => Dangling_Input_Signal,
       i_output_data_addr_reg(16) => Dangling_Input_Signal,
       i_output_data_addr_reg(17) => Dangling_Input_Signal,
       i_output_data_addr_reg(18) => Dangling_Input_Signal,
       i_output_data_addr_reg(19) => Dangling_Input_Signal,
       i_output_data_addr_reg(20) => Dangling_Input_Signal,
       i_output_data_addr_reg(21) => Dangling_Input_Signal,
       i_output_data_addr_reg(22) => Dangling_Input_Signal,
       i_output_data_addr_reg(23) => Dangling_Input_Signal,
       i_output_data_addr_reg(24) => Dangling_Input_Signal,
       i_output_data_addr_reg(25) => Dangling_Input_Signal,
       i_output_data_addr_reg(26) => Dangling_Input_Signal,
       i_output_data_addr_reg(27) => Dangling_Input_Signal,
       i_output_data_addr_reg(28) => Dangling_Input_Signal,
       i_output_data_addr_reg(29) => Dangling_Input_Signal,
       i_output_data_addr_reg(30) => Dangling_Input_Signal,
       i_output_data_addr_reg(31) => Dangling_Input_Signal,
       i_output_data_reg(0) => Dangling_Input_Signal,
       i_output_data_reg(1) => Dangling_Input_Signal,
       i_output_data_reg(2) => Dangling_Input_Signal,
       i_output_data_reg(3) => Dangling_Input_Signal,
       i_output_data_reg(4) => Dangling_Input_Signal,
       i_output_data_reg(5) => Dangling_Input_Signal,
       i_output_data_reg(6) => Dangling_Input_Signal,
       i_output_data_reg(7) => Dangling_Input_Signal,
       i_output_data_reg(8) => Dangling_Input_Signal,
       i_output_data_reg(9) => Dangling_Input_Signal,
       i_output_data_reg(10) => Dangling_Input_Signal,
       i_output_data_reg(11) => Dangling_Input_Signal,
       i_output_data_reg(12) => Dangling_Input_Signal,
       i_output_data_reg(13) => Dangling_Input_Signal,
       i_output_data_reg(14) => Dangling_Input_Signal,
       i_output_data_reg(15) => Dangling_Input_Signal,
       i_output_data_reg(16) => Dangling_Input_Signal,
       i_output_data_reg(17) => Dangling_Input_Signal,
       i_output_data_reg(18) => Dangling_Input_Signal,
       i_output_data_reg(19) => Dangling_Input_Signal,
       i_output_data_reg(20) => Dangling_Input_Signal,
       i_output_data_reg(21) => Dangling_Input_Signal,
       i_output_data_reg(22) => Dangling_Input_Signal,
       i_output_data_reg(23) => Dangling_Input_Signal,
       i_output_data_reg(24) => Dangling_Input_Signal,
       i_output_data_reg(25) => Dangling_Input_Signal,
       i_output_data_reg(26) => Dangling_Input_Signal,
       i_output_data_reg(27) => Dangling_Input_Signal,
       i_output_data_reg(28) => Dangling_Input_Signal,
       i_output_data_reg(29) => Dangling_Input_Signal,
       i_output_data_reg(30) => Dangling_Input_Signal,
       i_output_data_reg(31) => Dangling_Input_Signal,
       i_relu_control_reg(0) => Dangling_Input_Signal,
       i_relu_control_reg(1) => Dangling_Input_Signal,
       i_relu_control_reg(2) => Dangling_Input_Signal,
       i_relu_control_reg(3) => Dangling_Input_Signal,
       i_relu_control_reg(4) => Dangling_Input_Signal,
       i_relu_control_reg(5) => Dangling_Input_Signal,
       i_relu_control_reg(6) => Dangling_Input_Signal,
       i_relu_control_reg(7) => Dangling_Input_Signal,
       i_relu_control_reg(8) => Dangling_Input_Signal,
       i_relu_control_reg(9) => Dangling_Input_Signal,
       i_relu_control_reg(10) => Dangling_Input_Signal,
       i_relu_control_reg(11) => Dangling_Input_Signal,
       i_relu_control_reg(12) => Dangling_Input_Signal,
       i_relu_control_reg(13) => Dangling_Input_Signal,
       i_relu_control_reg(14) => Dangling_Input_Signal,
       i_relu_control_reg(15) => Dangling_Input_Signal,
       i_relu_control_reg(16) => Dangling_Input_Signal,
       i_relu_control_reg(17) => Dangling_Input_Signal,
       i_relu_control_reg(18) => Dangling_Input_Signal,
       i_relu_control_reg(19) => Dangling_Input_Signal,
       i_relu_control_reg(20) => Dangling_Input_Signal,
       i_relu_control_reg(21) => Dangling_Input_Signal,
       i_relu_control_reg(22) => Dangling_Input_Signal,
       i_relu_control_reg(23) => Dangling_Input_Signal,
       i_relu_control_reg(24) => Dangling_Input_Signal,
       i_relu_control_reg(25) => Dangling_Input_Signal,
       i_relu_control_reg(26) => Dangling_Input_Signal,
       i_relu_control_reg(27) => Dangling_Input_Signal,
       i_relu_control_reg(28) => Dangling_Input_Signal,
       i_relu_control_reg(29) => Dangling_Input_Signal,
       i_relu_control_reg(30) => Dangling_Input_Signal,
       i_relu_control_reg(31) => Dangling_Input_Signal,
       i_repeat_reg(0) => Dangling_Input_Signal,
       i_repeat_reg(1) => Dangling_Input_Signal,
       i_repeat_reg(2) => Dangling_Input_Signal,
       i_repeat_reg(3) => Dangling_Input_Signal,
       i_repeat_reg(4) => Dangling_Input_Signal,
       i_repeat_reg(5) => Dangling_Input_Signal,
       i_repeat_reg(6) => Dangling_Input_Signal,
       i_repeat_reg(7) => Dangling_Input_Signal,
       i_repeat_reg(8) => Dangling_Input_Signal,
       i_repeat_reg(9) => Dangling_Input_Signal,
       i_repeat_reg(10) => Dangling_Input_Signal,
       i_repeat_reg(11) => Dangling_Input_Signal,
       i_repeat_reg(12) => Dangling_Input_Signal,
       i_repeat_reg(13) => Dangling_Input_Signal,
       i_repeat_reg(14) => Dangling_Input_Signal,
       i_repeat_reg(15) => Dangling_Input_Signal,
       i_repeat_reg(16) => Dangling_Input_Signal,
       i_repeat_reg(17) => Dangling_Input_Signal,
       i_repeat_reg(18) => Dangling_Input_Signal,
       i_repeat_reg(19) => Dangling_Input_Signal,
       i_repeat_reg(20) => Dangling_Input_Signal,
       i_repeat_reg(21) => Dangling_Input_Signal,
       i_repeat_reg(22) => Dangling_Input_Signal,
       i_repeat_reg(23) => Dangling_Input_Signal,
       i_repeat_reg(24) => Dangling_Input_Signal,
       i_repeat_reg(25) => Dangling_Input_Signal,
       i_repeat_reg(26) => Dangling_Input_Signal,
       i_repeat_reg(27) => Dangling_Input_Signal,
       i_repeat_reg(28) => Dangling_Input_Signal,
       i_repeat_reg(29) => Dangling_Input_Signal,
       i_repeat_reg(30) => Dangling_Input_Signal,
       i_repeat_reg(31) => Dangling_Input_Signal,
       i_start_reg(0) => Dangling_Input_Signal,
       i_start_reg(1) => Dangling_Input_Signal,
       i_start_reg(2) => Dangling_Input_Signal,
       i_start_reg(3) => Dangling_Input_Signal,
       i_start_reg(4) => Dangling_Input_Signal,
       i_start_reg(5) => Dangling_Input_Signal,
       i_start_reg(6) => Dangling_Input_Signal,
       i_start_reg(7) => Dangling_Input_Signal,
       i_start_reg(8) => Dangling_Input_Signal,
       i_start_reg(9) => Dangling_Input_Signal,
       i_start_reg(10) => Dangling_Input_Signal,
       i_start_reg(11) => Dangling_Input_Signal,
       i_start_reg(12) => Dangling_Input_Signal,
       i_start_reg(13) => Dangling_Input_Signal,
       i_start_reg(14) => Dangling_Input_Signal,
       i_start_reg(15) => Dangling_Input_Signal,
       i_start_reg(16) => Dangling_Input_Signal,
       i_start_reg(17) => Dangling_Input_Signal,
       i_start_reg(18) => Dangling_Input_Signal,
       i_start_reg(19) => Dangling_Input_Signal,
       i_start_reg(20) => Dangling_Input_Signal,
       i_start_reg(21) => Dangling_Input_Signal,
       i_start_reg(22) => Dangling_Input_Signal,
       i_start_reg(23) => Dangling_Input_Signal,
       i_start_reg(24) => Dangling_Input_Signal,
       i_start_reg(25) => Dangling_Input_Signal,
       i_start_reg(26) => Dangling_Input_Signal,
       i_start_reg(27) => Dangling_Input_Signal,
       i_start_reg(28) => Dangling_Input_Signal,
       i_start_reg(29) => Dangling_Input_Signal,
       i_start_reg(30) => Dangling_Input_Signal,
       i_start_reg(31) => Dangling_Input_Signal,
       i_status_reg(0) => Dangling_Input_Signal,
       i_status_reg(1) => Dangling_Input_Signal,
       i_status_reg(2) => Dangling_Input_Signal,
       i_status_reg(3) => Dangling_Input_Signal,
       i_status_reg(4) => Dangling_Input_Signal,
       i_status_reg(5) => Dangling_Input_Signal,
       i_status_reg(6) => Dangling_Input_Signal,
       i_status_reg(7) => Dangling_Input_Signal,
       i_status_reg(8) => Dangling_Input_Signal,
       i_status_reg(9) => Dangling_Input_Signal,
       i_status_reg(10) => Dangling_Input_Signal,
       i_status_reg(11) => Dangling_Input_Signal,
       i_status_reg(12) => Dangling_Input_Signal,
       i_status_reg(13) => Dangling_Input_Signal,
       i_status_reg(14) => Dangling_Input_Signal,
       i_status_reg(15) => Dangling_Input_Signal,
       i_status_reg(16) => Dangling_Input_Signal,
       i_status_reg(17) => Dangling_Input_Signal,
       i_status_reg(18) => Dangling_Input_Signal,
       i_status_reg(19) => Dangling_Input_Signal,
       i_status_reg(20) => Dangling_Input_Signal,
       i_status_reg(21) => Dangling_Input_Signal,
       i_status_reg(22) => Dangling_Input_Signal,
       i_status_reg(23) => Dangling_Input_Signal,
       i_status_reg(24) => Dangling_Input_Signal,
       i_status_reg(25) => Dangling_Input_Signal,
       i_status_reg(26) => Dangling_Input_Signal,
       i_status_reg(27) => Dangling_Input_Signal,
       i_status_reg(28) => Dangling_Input_Signal,
       i_status_reg(29) => Dangling_Input_Signal,
       i_status_reg(30) => Dangling_Input_Signal,
       i_status_reg(31) => Dangling_Input_Signal,
       i_clk => Dangling_Input_Signal,
       i_reset_n => Dangling_Input_Signal
  );


---- Dangling input signal assignment ----

Dangling_Input_Signal <= DANGLING_INPUT_CONSTANT;

end arch;
